CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 80 1278 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
11
2 +V
167 150 156 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 950 287 0 17 19
10 12 11 10 9 8 7 6 18 2
1 1 1 1 0 0 1 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3536 0 0
2
5.89883e-315 0
0
7 Ground~
168 950 227 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89883e-315 0
0
7 Pulser~
4 71 233 0 10 12
0 19 20 4 4 0 0 5 5 2
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
5.89883e-315 0
0
6 74112~
219 383 269 0 7 32
0 5 17 4 17 5 21 16
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
3670 0 0
2
5.89883e-315 0
0
6 74LS48
188 874 371 0 14 29
0 13 15 16 17 22 23 6 7 8
9 10 11 12 24
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 695 141 0 3 22
0 3 15 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9323 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 489 132 0 3 22
0 17 16 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
317 0 0
2
5.89883e-315 0
0
6 74112~
219 775 263 0 7 32
0 5 14 4 14 5 25 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3108 0 0
2
5.89883e-315 0
0
6 74112~
219 569 267 0 7 32
0 5 3 4 3 5 26 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4299 0 0
2
5.89883e-315 0
0
6 74112~
219 197 269 0 7 32
0 5 5 4 5 5 27 17
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
9672 0 0
2
5.89883e-315 0
0
38
0 2 3 0 0 8192 0 0 10 29 0 3
536 234
536 231
545 231
0 1 3 0 0 4224 0 0 7 29 0 2
516 132
671 132
1 9 2 0 0 4224 0 3 2 0 0 2
950 235
950 245
4 0 4 0 0 4096 0 4 0 0 5 2
101 233
101 276
3 0 4 0 0 12288 0 4 0 0 35 5
95 224
101 224
101 276
163 276
163 323
5 0 5 0 0 4096 0 10 0 0 13 2
569 279
569 297
5 0 5 0 0 0 0 5 0 0 13 2
383 281
383 297
1 0 5 0 0 0 0 5 0 0 12 2
383 206
383 192
1 0 5 0 0 0 0 10 0 0 12 2
569 204
569 192
1 0 5 0 0 0 0 11 0 0 12 2
197 206
197 192
0 0 5 0 0 4096 0 0 0 12 13 2
287 192
287 297
0 1 5 0 0 4224 0 0 9 14 0 3
150 192
775 192
775 200
5 5 5 0 0 0 0 11 9 0 0 4
197 281
197 297
775 297
775 275
1 0 5 0 0 0 0 1 0 0 15 2
150 165
150 233
0 2 5 0 0 0 0 0 11 16 0 2
150 233
173 233
4 2 5 0 0 0 0 11 11 0 0 4
173 251
150 251
150 233
173 233
7 7 6 0 0 4224 0 6 2 0 0 3
906 335
965 335
965 323
8 6 7 0 0 4224 0 6 2 0 0 3
906 344
959 344
959 323
9 5 8 0 0 4224 0 6 2 0 0 3
906 353
953 353
953 323
10 4 9 0 0 4224 0 6 2 0 0 3
906 362
947 362
947 323
11 3 10 0 0 8320 0 6 2 0 0 3
906 371
941 371
941 323
12 2 11 0 0 8320 0 6 2 0 0 3
906 380
935 380
935 323
13 1 12 0 0 8320 0 6 2 0 0 3
906 389
929 389
929 323
7 1 13 0 0 8320 0 9 6 0 0 4
799 227
811 227
811 335
842 335
4 0 14 0 0 4096 0 9 0 0 26 3
751 245
720 245
720 227
2 3 14 0 0 8320 0 9 7 0 0 4
751 227
719 227
719 141
716 141
0 2 15 0 0 8320 0 0 6 28 0 3
657 231
657 344
842 344
7 2 15 0 0 0 0 10 7 0 0 4
593 231
658 231
658 150
671 150
4 3 3 0 0 0 0 10 8 0 0 6
545 249
536 249
536 231
516 231
516 132
510 132
3 0 4 0 0 8192 0 10 0 0 35 3
539 240
529 240
529 323
0 3 16 0 0 8320 0 0 6 32 0 3
461 233
461 353
842 353
7 2 16 0 0 0 0 5 8 0 0 4
407 233
461 233
461 141
465 141
4 0 17 0 0 4096 0 5 0 0 38 3
359 251
319 251
319 233
3 0 4 0 0 0 0 5 0 0 35 3
353 242
349 242
349 323
3 3 4 0 0 12416 0 11 9 0 0 6
167 242
163 242
163 323
737 323
737 236
745 236
0 4 17 0 0 8320 0 0 6 38 0 3
253 233
253 362
842 362
1 0 17 0 0 0 0 8 0 0 33 3
465 123
319 123
319 233
7 2 17 0 0 0 0 11 5 0 0 2
221 233
359 233
2
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
281 33 588 68
291 41 577 64
22 BINARY 4-BIT SYNCHRONO
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
566 33 756 68
576 41 745 64
13 US UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
